/* The Great Decider will take in keyboard input, 
who's player turn it is, and the players board

*/
module THE_GREAT_DECIDER ( 
	clock27 
	);
	input [1:0] clock27;
	
endmodule